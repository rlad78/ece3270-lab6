LIBRARY ieee;
USE ieee.std_logic_1164.all;


ENTITY bitpair_cl is
	PORT(clock, resetn, ivalid, iready: IN std_logic;
		  datain: IN std_logic_vector(31 downto 0);
		  oready, ovalid: OUT std_logic;
		  dataout: OUT std_logic_vector(31 downto 0));
END bitpair_cl;

ARCHITECTURE structure of bitpair_cl is
	

	BEGIN
		

END structure;
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
	
	
	
